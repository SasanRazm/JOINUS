.model jjmod jj(Rtype=1, Vg=2.71572mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=100uA)
.subckt jtl          1          2         3
R1                 3         4   8.34ohm
IR1   3   4   NOISE(5.274p 0.0 1.0p)
LPIN               1         5   0.354pH fcheck
LPR1               4         5   0.278pH fcheck
L2                 6         7   4.859pH fcheck
L3                 7         2   2.031pH fcheck
L1                 5         6   2.517pH fcheck
LP2                8         0   0.096pH fcheck
LP1                9         0   0.086pH fcheck
B2                 7         8  jjmod area=2.16
RS2                7         8   1.73ohm 
IRS2   7   8   NOISE(11.579p 0.0 1.0p)
B1                 6         9  jjmod area=2.16
RS1                6         9   1.73ohm 
IRS1   6   9   NOISE(11.579p 0.0 1.0p)
.ends
.subckt sink          1        10
R1                10        11   8.34ohm
IR1   10   11   NOISE(5.274p 0.0 1.0p)
R2                12         0   4.02ohm
IR2   12   0   NOISE(7.596p 0.0 1.0p)
LPIN               1        13   0.364pH fcheck
LPR1              11        13   0.265pH fcheck
L3                 9        12   5.307pH fcheck
L1                13         9   2.493pH fcheck
LP1                7         0   0.101pH fcheck
B1                 9         7  jjmod area=2.16
RS1                9         7   1.73ohm 
IRS1   9   7   NOISE(11.579p 0.0 1.0p)
.ends
.subckt SLTFF          1         14         15        17
L10               18        14   1.544pH fcheck
L11                8        15   2.350pH fcheck
LP7               19         0   0.190pH fcheck
L8                 7        18   3.097pH fcheck
L9                20         8   4.685pH fcheck
LP6               13         0   0.211pH fcheck
LPR2              21         7   0.520pH fcheck
L7                22         7   0.653pH fcheck
LP8               23        24   0.406pH fcheck
L12               25        22   0.003pH fcheck
L13               26        20   0.003pH fcheck
L5                23        22   3.146pH fcheck  
L6                20        23   3.214pH fcheck  
LP5               27         0   0.229pH fcheck
LP4               28         0   0.302pH fcheck
L2                29         9   1.019pH fcheck
L4                12         9   1.932pH fcheck  
L3                 9        30   1.851pH fcheck  
L1                31        29   2.369pH fcheck
LP1               32         0   0.130pH fcheck
LPR1              33        31   0.247pH fcheck
LPDIN              1        31   0.218pH fcheck
RD                24         0   2.00ohm           
IRD   24   0   NOISE(10.769p 0.0 1.0p)
R2                17        21  16.67ohm
IR2   17   21   NOISE(3.73p 0.0 1.0p)
R1                17        33   8.34ohm
IR1   17   33   NOISE(5.274p 0.0 1.0p)
B7                 8        19  jjmod area=2.18
RS7                8        19   1.71ohm 
IRS7   8   19   NOISE(11.646p 0.0 1.0p)
B6                18        13  jjmod area=2.18
RS6               18        13   1.71ohm 
IRS6   18   13   NOISE(11.646p 0.0 1.0p)
B5                26        27  jjmod area=1.96
RS5               26        27   1.90ohm 
IRS5   26   27   NOISE(11.049p 0.0 1.0p)
B3                26        12  jjmod area=1.32      
RS3               26        12   2.83ohm 
IRS3   26   12   NOISE(9.053p 0.0 1.0p)
B2                25        30  jjmod area=1.84      
RS2               25        30   2.03ohm 
IRS2   25   30   NOISE(10.689p 0.0 1.0p)
B4                25        28  jjmod area=1.10
RS4               25        28   3.39ohm 
IRS4   25   28   NOISE(8.272p 0.0 1.0p)
B1                29        32  jjmod area=2.18
RS1               29        32   1.71ohm 
IRS1   29   32   NOISE(11.646p 0.0 1.0p)
K1                L5        L6   -0.14
.ends
Vclk              36          0  PULSE(0.0mV  1.034mV   0ps   1.0ps   1.0ps   1.0ps   30.0ps)
XI0               jtl         36         34         37
XI1               jtl         34         35         37
XI4             SLTFF         35         31         29         37
XI6               jtl         29         26         37
XI2              sink         26         37
XI5               jtl         31         10         37
XI7             SLTFF         10         50         51         37
XI14               jtl         51         52         37
XI3              sink         52         37
XI8               jtl         50         53         37
XI9             SLTFF         53         54         55         37
XI10               jtl         55         56         37
XI11              sink         56         37
XI12              sink         54         37
V1                37         0  PWL(0ps 0mv 10ps 2.5mv)
.tran 0.5PS 5nS 10PS 0.1PS
.file OUTCNT.DAT
.print Devv XI1_B2
.print Devv XI2_B1
.print Devv XI3_B1
.print Devv XI11_B1
