*** Example for the I-V charascteristic and the Shapiro step with microwave pumping 
*** for a damped Josephson junction.

*JSIM model
.model jjmod jj(Rtype=1, Vg=2.8mV, Cap=0.218pF, R0=200ohm, Rn=17ohm, Icrit=0.1mA)

*** netlist file ***
**** **** **** **** **** **** **** ****+
*** Lib : Example1
*** Cell: JJIV
*** View: Schematic
*** Jan 2019
**** **** **** **** **** **** **** ****

*** ptl_2ohm
.subckt ptl_2ohm          2          3
***       din      dout
C1                 2         0   0.168pF
L1                 2         3   0.665pH fcheck
.ends

*** top cell: JJ210
B8                1        2   jjmod area=2.20
RS8               1        2   1.70ohm *SHUNT=3.73
XI1        ptl_2ohm  1        3   
Rsource           3        0   1000ohm
Rsource2	  2       0   1ohm
I0                0        1   PWL(0ps 0mA 100ps 1mA)


*** jsim input file ***
.tran 0.01ps 150PS 100PS 0.1PS
.FILE OUT.DAT
.PRINT DEVI Rsource2
.PRINT nodev 1 0